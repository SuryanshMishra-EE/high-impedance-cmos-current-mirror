* C:\Users\Suryansh Mishra\Documents\Ltspice_schematics\schematic_output_impedance.asc
M1 N003 N003 N007 N007 CMOSN l=180nm w=360nm
M2 N004 N004 N007 N007 CMOSN l=180nm w=360nm
M3 N007 N004 0 0 CMOSN l=180nm w=360nm
M4 vdd N004 N008 N008 CMOSN l=180nm w=360nm
M5 N004 N004 N008 N008 CMOSN l=180nm w=360nm
M6 N008 N004 0 0 CMOSN l=180nm w=360nm
I1 0 N003 40µ
I2 0 N004 40µ
I3 0 N004 40µ
M7 N012 N011 N013 N013 CMOSN l=360nm w=204nm
M8 N013 N011 0 0 CMOSN l=360nm w=568nm
M9 vdd N012 N014 N014 CMOSN l=360nm w=364nm
M10 N011 N011 N014 N014 CMOSN l=360nm w=204nm
M11 N014 N011 0 0 CMOSN l=360nm w=568nm
M12 N010 N009 N012 N010 CMOSP l=360nm w=403nm
M13 N010 N009 N011 N010 CMOSP l=360nm w=403nm
V2 N010 0 1.8
V3 N009 0 2.1
I4 0 N013 5µ
Vbias vdd 0 1.8
M15 N002 N001 N005 N005 CMOSN l=180nm w=360nm
M16 N005 N001 0 0 CMOSN l=180nm w=360nm
M17 N001 N001 N006 N006 CMOSN l=180nm w=360nm
M18 vdd N002 N006 N006 CMOSN l=180nm w=360nm
I6 0 N005 40µ
I7 0 N002 40µ
I8 0 N001 40µ
M19 N006 N001 0 0 CMOSN l=180nm w=360nm
.model NMOS NMOS
.model PMOS PMOS
.lib C:\Users\Suryansh Mishra\AppData\Local\LTspice\lib\cmp\standard.mos
.INCLUDE tsmc018.lib
.INCLUDE tsmc018.lib
.INCLUDE tsmc018.lib
.dc Vbias 0.501 1.8 0.25
.backanno
.end
